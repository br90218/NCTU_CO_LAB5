//Subject:		CO project 5 - Sign extend
//--------------------------------------------------------------------------------
//Version:		1
//--------------------------------------------------------------------------------
//Writer:		0210022 鍾承佑, 0210029 鄧仰哲
//----------------------------------------------
//Date:
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );

//I/O ports
input	[16-1:0]	data_i;
output	[32-1:0]	data_o;

//Internal Signals
reg		[32-1:0]	data_o;

//Sign extended
always@ (data_i) begin
	if (data_i[15]==1'b1)
		data_o[31 -: 16]=16'b1111111111111111;
	else
		data_o[31 -: 16]=16'b0;

	data_o[15 -: 16]=data_i;
end

endmodule