//Subject:		CO project 5 - Shift_Left_Two_32
//--------------------------------------------------------------------------------
//Version:		1
//--------------------------------------------------------------------------------
//Writer:		0210022 鍾承佑, 0210029 鄧仰哲
//----------------------------------------------
//Date:
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Shift_Left_Two_32(
    data_i,
    data_o
    );

//I/O ports
input	[32-1:0]	data_i;
output	[32-1:0]	data_o;

//shift left 2
assign data_o[32-1 -: 30] = data_i[29:0];
assign data_o[1:0] = 2'b00;

endmodule